module memory_led (
    input led
    output addr
    output addr_side
);

always @ (negedge clk) begin
    
end

endmodule